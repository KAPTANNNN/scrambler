//module scrambler (
 //   input clk,
 //   input reset,
 //   input serial_input,
 //   output reg [7:0] scrambled_output // Define width of the output explicitly
//);
   // wire [14:0] lfsr_out;

   // lfsr lfsr_inst (
     //   .clk(clk),
      //  .reset(reset),
       // .lfsr_out(lfsr_out)
   // );

   // always @(posedge clk or posedge reset) begin
       // if (reset)
        //    scrambled_output <= 8'b0;
        //else
        //    scrambled_output <= serial_input ^ lfsr_out[14]; // Scramble the input bit
    //end//
//endmodule
